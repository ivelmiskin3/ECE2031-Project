LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

LIBRARY WORK;

ENTITY SLOW_SRAM IS
  PORT (
    IO_WRITE : IN STD_LOGIC;
    SRAM_ADLOW_EN : IN STD_LOGIC;
    SRAM_ADHI_EN : IN STD_LOGIC;
    SRAM_DATA_EN : IN STD_LOGIC;
    SRAM_CTRL_EN : IN STD_LOGIC;
    IO_DATA : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    SRAM_DQ : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    SRAM_CE_N : OUT STD_LOGIC;
    SRAM_WE_N : OUT STD_LOGIC;
    SRAM_OE_N : OUT STD_LOGIC;
    SRAM_UB_N : OUT STD_LOGIC;
    SRAM_LB_N : OUT STD_LOGIC;
    SRAM_ADDR : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END SLOW_SRAM;

ARCHITECTURE BDF_TYPE OF SLOW_SRAM IS

  COMPONENT LPM_BUSTRI_OE0
    PORT (
      enabledt : IN STD_LOGIC;
      data : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
      tridata : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0)
    );
  END COMPONENT;

  COMPONENT LPM_FF0
    PORT (
      clock : IN STD_LOGIC;
      data : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
      q : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
    );
  END COMPONENT;

  COMPONENT LPM_FF1
    PORT (
      clock : IN STD_LOGIC;
      data : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      q : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
    );
  END COMPONENT;

  SIGNAL SRAM_ADDR_ALTERA : STD_LOGIC_VECTOR(17 DOWNTO 0);
  SIGNAL SRAM_CTRL : STD_LOGIC_VECTOR(2 DOWNTO 0);
  SIGNAL SRAM_IO_DATA : STD_LOGIC_VECTOR(15 DOWNTO 0);

BEGIN
  SRAM_CE_N <= '0';
  SRAM_UB_N <= '0';
  SRAM_LB_N <= '0';

  OUTPUT_BUS : LPM_BUSTRI_OE0
  PORT MAP(
    enabledt => SRAM_CTRL(2),
    data => SRAM_IO_DATA,
    tridata => SRAM_DQ
  );

  INPUT_BUS : LPM_BUSTRI_OE0
  PORT MAP(
    enabledt => NOT(IO_WRITE) AND SRAM_DATA_EN,
    data => SRAM_DQ,
    tridata => IO_DATA
  );

  ADDR_LB : LPM_FF0
  PORT MAP(
    clock => IO_WRITE AND SRAM_ADLOW_EN,
    data => IO_DATA,
    q => SRAM_ADDR_ALTERA(15 DOWNTO 0)
  );

  IO_REGISTER : LPM_FF0
  PORT MAP(
    clock => SRAM_DATA_EN AND IO_WRITE,
    data => IO_DATA,
    q => SRAM_IO_DATA
  );

  ADDR_UB : LPM_FF1
  PORT MAP(
    clock => IO_WRITE AND SRAM_ADHI_EN,
    data => IO_DATA(1 DOWNTO 0),
    q => SRAM_ADDR_ALTERA(17 DOWNTO 16)
  );

  CONTROL : LPM_FF1
  PORT MAP(
    clock => IO_WRITE AND SRAM_CTRL_EN,
    data => IO_DATA(2 DOWNTO 0),
    q => SRAM_CTRL
  );

  SRAM_WE_N <= SRAM_CTRL(1);
  SRAM_OE_N <= SRAM_CTRL(0);
  SRAM_ADDR <= SRAM_ADDR_ALTERA;

END BDF_TYPE;