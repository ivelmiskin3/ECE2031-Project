LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
use ieee.numeric_std.all;

LIBRARY work;

ENTITY addressimplementation IS
  PORT (
    IO_WRITE : IN STD_LOGIC;
    SRAM_SET_UPPER : IN STD_LOGIC;
    SRAM_SET_LOWER : IN STD_LOGIC;
    SRAM_DATA : IN STD_LOGIC;
    SRAM_INC_DATA : IN STD_LOGIC;
    IO_DATA : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    SRAM_CE_N : OUT STD_LOGIC;
    SRAM_WE_N : OUT STD_LOGIC;
    SRAM_OE_N : OUT STD_LOGIC;
    SRAM_UB_N : OUT STD_LOGIC;
    SRAM_LB_N : OUT STD_LOGIC;
    SRAM_ADDR : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END addressimplementation;

ARCHITECTURE bdf_type OF addressimplementation IS
  SIGNAL SRAM_ADDR_ALTERA_SYNTHESIZED : STD_LOGIC_VECTOR(17 DOWNTO 0);
  SIGNAL UPPER_ENABLE : boolean;
  SIGNAL LOWER_ENABLE : boolean;
  SIGNAL WRITE_ENABLE : boolean;
  SIGNAL READ_ENABLE : boolean;
--  SIGNAL INCREMENT_ADDRESS : boolean;
BEGIN
  -- Default SRAM Control Signals
  SRAM_CE_N <= '0';
  SRAM_UB_N <= '0';
  SRAM_LB_N <= '0';
  SRAM_ADDR <= SRAM_ADDR_ALTERA_SYNTHESIZED;
  
  -- Actions
  UPPER_ENABLE <= SRAM_SET_UPPER = '1' AND IO_WRITE = '1';
  LOWER_ENABLE <= SRAM_SET_LOWER = '1' AND IO_WRITE = '1';
  WRITE_ENABLE <= (SRAM_DATA = '1' OR SRAM_INC_DATA = '1') AND IO_WRITE = '1';
  READ_ENABLE <= (SRAM_DATA = '1' OR SRAM_INC_DATA = '1') AND IO_WRITE = '0';
  
  PROCESS (UPPER_ENABLE, LOWER_ENABLE, WRITE_ENABLE, READ_ENABLE)
  BEGIN
	-- SET UPPER
	IF UPPER_ENABLE THEN
		SRAM_ADDR_ALTERA_SYNTHESIZED(17 DOWNTO 16) <= IO_DATA(1 DOWNTO 0);
	END IF;
	
	-- SET LOWER
	IF LOWER_ENABLE THEN
		SRAM_ADDR_ALTERA_SYNTHESIZED(15 DOWNTO 0) <= IO_DATA(15 DOWNTO 0);
	END IF;
	
	-- READ OR WRITE
	IF WRITE_ENABLE AND NOT READ_ENABLE THEN
		SRAM_WE_N <= '0';
	ELSIF READ_ENABLE AND NOT WRITE_ENABLE THEN
		SRAM_OE_N <= '0';
	ELSE
		SRAM_WE_N <= '1';
		SRAM_OE_N <= '1';
	END IF;
	
	-- INCREMENT
--	IF (SRAM_INC_DATA = '1') THEN
--		INCREMENT_ADDRESS <= true;
--	ELSIF (INCREMENT_ADDRESS AND SRAM_INC_DATA = '0') THEN
--		INCREMENT_ADDRESS <= false;
--		SRAM_ADDR_VHDL_SYNTHESIZED <= std_logic_vector(unsigned(SRAM_ADDR_VHDL_SYNTHESIZED) + 1);
--	END IF;
  END PROCESS;
END bdf_type;